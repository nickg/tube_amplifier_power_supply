library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package tubepsu_addresses_pkg is



end package tubepsu_addresses_pkg;
